`define s_IO_READ ($fell (framen) && (cxben[3:0] == 4'b0010))
