`define s_IO_READ         ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_IO_WRITE        ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_MEM_READ        ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_MEM_WRITE       ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_CONFIG_READ     ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_CONFIG_WRITE    ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_DUAL_ADDR_CYCLE ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_MEM_READ_LINE   ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_MEM_WRITE_INV   ($fell (framen) && (cxben[3:0] == 4'b0010))
`define s_BUS_IDLE        ($fell (framen) && (cxben[3:0] == 4'b0010))
